library verilog;
use verilog.vl_types.all;
entity Rtype_testbench2 is
end Rtype_testbench2;
