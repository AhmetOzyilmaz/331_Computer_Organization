library verilog;
use verilog.vl_types.all;
entity Rtype_testbench is
end Rtype_testbench;
