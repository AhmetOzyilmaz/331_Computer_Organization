library verilog;
use verilog.vl_types.all;
entity project01 is
    port(
        R               : out    vl_logic_vector(4 downto 0);
        A               : in     vl_logic_vector(4 downto 0);
        B               : in     vl_logic_vector(4 downto 0);
        S               : in     vl_logic_vector(1 downto 0)
    );
end project01;
