module mips_testbench ();

reg [31:0] instruction_set;
wire result;

initial begin
instruction_set = 32'b00000010000100101000000100000; #10;
//....continue for all instruction types.... must be least 9 control

end






endmodule