module mips_core(instruction, result);

input [31:0] instruction;
output [31:0] result;









endmodule