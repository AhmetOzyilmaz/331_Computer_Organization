library verilog;
use verilog.vl_types.all;
entity FivebitAnd_Testbench is
end FivebitAnd_Testbench;
