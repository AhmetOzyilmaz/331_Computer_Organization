library verilog;
use verilog.vl_types.all;
entity project01_Testbench is
end project01_Testbench;
